 `include "define.v"
module ysyx_25060170_top (
    input clk,
    input rst
);


endmodule

